module sim_pc_irom ();
  reg clk;
    
endmodule