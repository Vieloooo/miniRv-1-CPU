module top (
    input clk,
    input halt
);

    
endmodule